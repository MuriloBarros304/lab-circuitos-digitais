library verilog;
use verilog.vl_types.all;
entity mux8b_vlg_vec_tst is
end mux8b_vlg_vec_tst;
