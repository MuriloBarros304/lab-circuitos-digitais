library verilog;
use verilog.vl_types.all;
entity regFlipflop_vlg_vec_tst is
end regFlipflop_vlg_vec_tst;
