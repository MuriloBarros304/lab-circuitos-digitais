library verilog;
use verilog.vl_types.all;
entity calc_vlg_vec_tst is
end calc_vlg_vec_tst;
