library verilog;
use verilog.vl_types.all;
entity decrementador_vlg_vec_tst is
end decrementador_vlg_vec_tst;
