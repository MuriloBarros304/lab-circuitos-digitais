library verilog;
use verilog.vl_types.all;
entity circuito_vlg_vec_tst is
end circuito_vlg_vec_tst;
