library verilog;
use verilog.vl_types.all;
entity mux2x1pl_vlg_vec_tst is
end mux2x1pl_vlg_vec_tst;
