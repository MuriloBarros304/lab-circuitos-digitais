library verilog;
use verilog.vl_types.all;
entity mux4x1pl_vlg_vec_tst is
end mux4x1pl_vlg_vec_tst;
