library verilog;
use verilog.vl_types.all;
entity d7segcomp_vlg_vec_tst is
end d7segcomp_vlg_vec_tst;
