library verilog;
use verilog.vl_types.all;
entity d7seg_vlg_vec_tst is
end d7seg_vlg_vec_tst;
