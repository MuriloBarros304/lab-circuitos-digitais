library verilog;
use verilog.vl_types.all;
entity regLatch_vlg_vec_tst is
end regLatch_vlg_vec_tst;
