library verilog;
use verilog.vl_types.all;
entity latchd_vlg_vec_tst is
end latchd_vlg_vec_tst;
